
library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM IS
   generic (
		dataWidth: natural := 32;
		addrWidth: natural := 32;
		memoryAddrWidth:  natural := 6 
	 );   -- 64 posicoes de 32 bits cada
   port ( 
		clk: IN  STD_LOGIC;
		Endereco: IN  STD_LOGIC_VECTOR (addrWidth-1 DOWNTO 0);
		Dado: OUT STD_LOGIC_VECTOR (dataWidth-1 DOWNTO 0) 
	);
end entity;

architecture assincrona OF ROM IS
  type blocoMemoria IS ARRAY(0 TO 2**memoryAddrWidth - 1) OF std_logic_vector(dataWidth-1 DOWNTO 0);
  
  signal memROM: blocoMemoria;
  attribute ram_init_file : string;
  attribute ram_init_file of memROM:
  signal is "MIPS_Intermediaria.mif";

   signal EnderecoLocal : std_logic_vector(memoryAddrWidth-1 downto 0);

begin
  EnderecoLocal <= Endereco(memoryAddrWidth+1 downto 2);
  Dado <= memROM (to_integer(unsigned(EnderecoLocal)));
end architecture;