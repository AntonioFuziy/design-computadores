library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Decoder is

  port   (
    -- Input ports
	 OPCODE: in std_logic_vector(3 downto 0);
	 OUTPUT: out std_logic_vector(10 downto 0)
  );
end entity;


architecture arch_name of Decoder is
  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101"; 
  constant JMP  : std_logic_vector(3 downto 0) := "0110"; 
  constant JEQ  : std_logic_vector(3 downto 0) := "0111"; 
  constant CEQ  : std_logic_vector(3 downto 0) := "1000"; 
  constant JSR  : std_logic_vector(3 downto 0) := "1001"; 
  constant RET  : std_logic_vector(3 downto 0) := "1010"; 
begin
	OUTPUT <= "00000011001" when OPCODE = LDA else
				 "00000010101" when OPCODE = SOMA else
				 "00000010001" when OPCODE = SUB else
				 "00000111000" when OPCODE = LDI else
				 "10000000000" when OPCODE = STA else
				 "01000000000" when OPCODE = JMP else
				 "01001000010" when OPCODE = JEQ else
				 "00000001111" when OPCODE = CEQ else
				 "11010000000" when OPCODE = JSR else
				 "01100000000" when OPCODE = RET else
				 "00000000000";
end architecture;